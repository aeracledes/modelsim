module pcoder(D3,D2,D1,D0,Y1,Y0,Z);

input D3,D2,D1,D0;
output reg Y1,Y0,Z;

always @(*)
	case ({D3,D2,D1,D0})
		4'b0000: {Y1,Y0,Z} = 3'b001;
		4'b0001: {Y1,Y0,Z} = 3'b000;
		4'b0010: {Y1,Y0,Z} = 3'b010;
		4'b0011: {Y1,Y0,Z} = 3'b010;
		4'b0100: {Y1,Y0,Z} = 3'b100;	
		4'b0101: {Y1,Y0,Z} = 3'b100;
		4'b0110: {Y1,Y0,Z} = 3'b100;
		4'b0111: {Y1,Y0,Z} = 3'b100;
		4'b1000: {Y1,Y0,Z} = 3'b110;
		4'b1001: {Y1,Y0,Z} = 3'b110;
		4'b1010: {Y1,Y0,Z} = 3'b110;
		4'b1011: {Y1,Y0,Z} = 3'b110;
		4'b1100: {Y1,Y0,Z} = 3'b110;
		4'b1101: {Y1,Y0,Z} = 3'b110;
		4'b1110: {Y1,Y0,Z} = 3'b110;
		4'b1111: {Y1,Y0,Z} = 3'b110;
	endcase
endmodule
	

